library verilog;
use verilog.vl_types.all;
entity image_vlg_vec_tst is
end image_vlg_vec_tst;
