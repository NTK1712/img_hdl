library verilog;
use verilog.vl_types.all;
entity sobel_vlg_vec_tst is
end sobel_vlg_vec_tst;
