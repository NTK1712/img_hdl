library verilog;
use verilog.vl_types.all;
entity test_gray is
end test_gray;
