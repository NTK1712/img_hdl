library verilog;
use verilog.vl_types.all;
entity test_image is
end test_image;
