library verilog;
use verilog.vl_types.all;
entity B_vlg_vec_tst is
end B_vlg_vec_tst;
