library verilog;
use verilog.vl_types.all;
entity test_sobel is
end test_sobel;
