library verilog;
use verilog.vl_types.all;
entity test_blur is
end test_blur;
